// syncfifo_w9d128_aclr_showahead.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module syncfifo_w9d128_aclr_showahead (
		input  wire [8:0] data,  //  fifo_input.datain
		input  wire       wrreq, //            .wrreq
		input  wire       rdreq, //            .rdreq
		input  wire       clock, //            .clk
		input  wire       aclr,  //            .aclr
		output wire [8:0] q,     // fifo_output.dataout
		output wire [6:0] usedw, //            .usedw
		output wire       full,  //            .full
		output wire       empty  //            .empty
	);

	syncfifo_w9d128_aclr_showahead_fifo_191_sqyurki fifo_0 (
		.data  (data),  //  fifo_input.datain
		.wrreq (wrreq), //            .wrreq
		.rdreq (rdreq), //            .rdreq
		.clock (clock), //            .clk
		.aclr  (aclr),  //            .aclr
		.q     (q),     // fifo_output.dataout
		.usedw (usedw), //            .usedw
		.full  (full),  //            .full
		.empty (empty)  //            .empty
	);

endmodule
